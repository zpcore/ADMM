LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;

library ADMM_lib;
use ADMM_lib.ADMM_pkg.all;
 
ENTITY ADMM_TOP_tb IS
END ADMM_TOP_tb;
 
ARCHITECTURE behavior OF ADMM_TOP_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
component ADMM_TOP is
	Port ( 
		CLK : in  STD_LOGIC;
		RST : in  STD_LOGIC;
		NumBRAM : in STD_LOGIC_VECTOR(31 downto 0);
		ADDRBRAM : in STD_LOGIC_VECTOR(31 downto 0);
		WRBRAM : in STD_LOGIC;
		MATData : in STD_LOGIC_VECTOR(31 downto 0);
		ConfigSTATE : in state_type;
--		START : in STD_LOGIC;--start computation signal, after BRAMInit state
		RHO : in STD_LOGIC_VECTOR(31 downto 0);
		ALPHA : in STD_LOGIC_VECTOR(31 downto 0);
		ONEMINUSALPHA : in STD_LOGIC_VECTOR(31 downto 0);
		U : out Mby32_type;
		STATE_RD : out STD_LOGIC;
		X : in STD_LOGIC_VECTOR(31 downto 0);--signal from sensor, serial input(x0,x1,...xN)
--below signal for simulation
		BOX : in STD_LOGIC_VECTOR(31 downto 0);
		BOX_REQUEST : out STD_LOGIC;
		QR : in STD_LOGIC_VECTOR(31 downto 0);
		NEW_QR_RDY : in STD_LOGIC
);
end component;

--Inputs
signal CLK : std_logic := '0';
signal RST : std_logic := '0';
signal NumBRAM : std_logic_vector(31 downto 0) := (others=>'0');
signal ADDRBRAM : std_logic_vector(31 downto 0) := (others=>'0');
signal WRBRAM : std_logic := '0';
signal MATData : std_logic_vector(31 downto 0) := (others=> '0');
signal ConfigSTATE : state_type := idle;
--signal START : std_logic := '0';
signal RHO : std_logic_vector(31 downto 0) := (others=>'0');
signal ALPHA : std_logic_vector(31 downto 0) := (others=>'0');
signal ONEMINUSALPHA : std_logic_vector(31 downto 0) := (others=>'0');
signal BOX : std_logic_vector(31 downto 0) := (others=>'0');
signal BOX_REQUEST : std_logic := '0';
signal QR : std_logic_vector(31 downto 0) := (others=>'0');
signal NEW_QR_RDY : std_logic := '0';
signal X : std_logic_vector(31 downto 0):=(others=>'0');
signal STATE_RD : std_logic:='0';

--Outputs
signal U : Mby32_type;

-- Clock period definitions
constant CLK_period : time := 10 ns;
 
BEGIN
 
-- Instantiate the Unit Under Test (UUT)
uut: ADMM_TOP PORT MAP (
	CLK =>CLK,
	RST =>RST,
	NumBRAM =>NumBRAM,
	ADDRBRAM =>ADDRBRAM,
	WRBRAM =>WRBRAM,
	MATData =>MATData,
	ConfigSTATE =>ConfigSTATE,
	RHO =>RHO,
	ALPHA =>ALPHA,
	ONEMINUSALPHA =>ONEMINUSALPHA,
	U =>U,
	STATE_RD => STATE_RD,
	X => X,
	--below signal for simulation
	BOX =>BOX,
	BOX_REQUEST =>BOX_REQUEST,
	QR =>QR,
	NEW_QR_RDY =>NEW_QR_RDY
	);

   -- Clock process definitions
CLK_process :process
begin
	CLK <= '0';
	wait for CLK_period/2;
	CLK <= '1';
	wait for CLK_period/2;
end process;

boxQR: process
begin		
	BOX <= x"425c0000";--55
	X <= x"3F800000";
	wait;
end process;

   -- Stimulus process
stim_proc: process
begin		
	-- hold reset state for 100 ns.
	RST <= '1';
	wait for 105.1 ns;	
  	RST <= '0';
	ALPHA <= x"3FC00000";--1.5
	ONEMINUSALPHA <= x"BF000000";-- -0.5
	RHO <= x"3F666666";--0.9
	QR <= x"00000000";
	wait for CLK_period*10;
	ConfigSTATE <= BRAM_init;

	wait for CLK_period;
	WRBRAM <= '1';
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(0,ADDRBRAM'length));
	MATData <= x"4085f20e";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(0,ADDRBRAM'length));
	MATData <= x"3fe025a0";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(0,ADDRBRAM'length));
	MATData <= x"410fc3a8";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(0,ADDRBRAM'length));
	MATData <= x"40ee0af0";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(1,ADDRBRAM'length));
	MATData <= x"406a8bcb";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(1,ADDRBRAM'length));
	MATData <= x"41149a27";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(1,ADDRBRAM'length));
	MATData <= x"40889e70";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(1,ADDRBRAM'length));
	MATData <= x"00000000";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2,ADDRBRAM'length));
	MATData <= x"4102803a";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2,ADDRBRAM'length));
	MATData <= x"3fcad588";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2,ADDRBRAM'length));
	MATData <= x"40daddd9";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2,ADDRBRAM'length));
	MATData <= x"410acfcb";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(3,ADDRBRAM'length));
	MATData <= x"40d01c56";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(3,ADDRBRAM'length));
	MATData <= x"410bf2d8";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(3,ADDRBRAM'length));
	MATData <= x"40b72f2c";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(3,ADDRBRAM'length));
	MATData <= x"00000000";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(4,ADDRBRAM'length));
	MATData <= x"40be09ae";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(4,ADDRBRAM'length));
	MATData <= x"40d03f71";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(4,ADDRBRAM'length));
	MATData <= x"4107d55a";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(4,ADDRBRAM'length));
	MATData <= x"3faf26ee";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(5,ADDRBRAM'length));
	MATData <= x"40ea641a";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(5,ADDRBRAM'length));
	MATData <= x"40961dd7";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(5,ADDRBRAM'length));
	MATData <= x"40ee26af";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(5,ADDRBRAM'length));
	MATData <= x"00000000";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(6,ADDRBRAM'length));
	MATData <= x"3fd1e298";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(6,ADDRBRAM'length));
	MATData <= x"40db2186";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(6,ADDRBRAM'length));
	MATData <= x"4108aa71";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(6,ADDRBRAM'length));
	MATData <= x"40b7f4a4";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(7,ADDRBRAM'length));
	MATData <= x"3f808d33";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(7,ADDRBRAM'length));
	MATData <= x"3fe00bbe";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(7,ADDRBRAM'length));
	MATData <= x"3f81acc1";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(7,ADDRBRAM'length));
	MATData <= x"00000000";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(8,ADDRBRAM'length));
	MATData <= x"407f5fa8";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(8,ADDRBRAM'length));
	MATData <= x"40c5ef2d";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(8,ADDRBRAM'length));
	MATData <= x"403e9138";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(8,ADDRBRAM'length));
	MATData <= x"40e5f33e";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(9,ADDRBRAM'length));
	MATData <= x"40efa902";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(9,ADDRBRAM'length));
	MATData <= x"4113d582";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(9,ADDRBRAM'length));
	MATData <= x"41112367";

	wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(9,ADDRBRAM'length));
	MATData <= x"00000000";
--------write vector
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2016,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2016,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2016,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2016,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(0, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2017,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(1, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2017,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(2, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2017,ADDRBRAM'length));
	MATData <= x"3f800000";
wait for CLK_period;
	NumBRAM <= std_logic_vector(to_unsigned(3, NumBRAM'length));
	ADDRBRAM <= std_logic_vector(to_unsigned(2017,ADDRBRAM'length));
	MATData <= x"3f800000";
-------write vector

	wait for CLK_period;
	WRBRAM <= '0';
	ConfigSTATE <= idle;	
	wait for CLK_period;
	ConfigSTATE <= QR_init;
	
	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fe5a535";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e3dc4b3";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fbb3879";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3eb15f94";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f9ddf62";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd88f3b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ff85f2f";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f9bb481";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f0674e6";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f914c4d";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fa74e8b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e330255";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fafe9be";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3eaf6e5a";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f720fdb";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f91c419";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f8c8e54";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f1bbd49";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ff760bf";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ff4dce9";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f5c7a94";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ed44bbc";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3feb82cf";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e062a41";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd105cb";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f11affe";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fe723f2";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e6dbc0b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ffe6f1a";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fb3d4c5";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f8d0444";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd8ae1b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ebffd01";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f333b3c";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ff48728";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e0f67a3";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f59302e";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f2148fb";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e8498e2";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fa1ecd9";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fcf3c1b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f9d70f8";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fa299a0";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f56680d";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f9f4cd5";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3eeb9aaa";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ea93b6b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ed3394d";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f47eadf";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f710d43";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f99c982";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f56e543";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f427764";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fb39b85";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e39c14b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ff3cadc";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e678a30";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f0c5f9e";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e8a5377";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd91f7e";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f248abd";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3dcda390";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fb53798";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f7373ed";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd49592";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f9c3292";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd4fd1a";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f8e086b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f4787b6";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f26420e";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3edb7fb8";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3efe9d54";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ebd090a";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e2daaf1";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fe3cdc3";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f37d48d";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f85d101";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fd85bf5";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fb8cddb";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f2a5ba1";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fc3a7da";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f71d3d8";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3e7a5b30";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fe9631b";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fc69ff0";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ee28e04";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f489cf1";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f7e694c";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3ef8b63f";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f396f17";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f8b49ab";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3dcfee84";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fc866dd";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3faa4ead";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fbb306a";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fee6cfd";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f18a172";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f783507";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3f71a3e3";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	wait for 2*CLK_period;
	NEW_QR_RDY <= '1';
	QR <= x"3fb63152";
	wait for CLK_period;
	NEW_QR_RDY <= '0';

	ConfigSTATE <= running;


	wait;
end process;



END;
